
module rkv_watchdog_tb;

    cmsdk_apb_watchdog dut();
    
endmodule
