`ifndef RKV_WATCHDOG_SEQ_LIB_SVH
`define RKV_WATCHDOG_SEQ_LIB_SVH

    `include"rkv_watchdog_base_virtual_sequence.sv"
    `include"rkv_watchdog_integration_virt_seq.sv"
    `include"rkv_watchdog_apbacc_virt_seq.sv"
    `include"rkv_watchdog_regacc_virt_seq.sv"


`endif // RKV_WATCHDOG_SEQ_LIB_SVH
