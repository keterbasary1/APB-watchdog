`ifndef RKV_WATCHDOG_CONFIG_SV
`define RKV_WATCHDOG_CONFIG_SV

class rkv_watchdog_config extends uvm_object;

    function new(string name = "rkv_watchdog_config");
        super.new(name);
    endfunction
    
endclass

`endif